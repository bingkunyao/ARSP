 
module altaccumulate_ref (cin, data, add_sub, clock, sload, clken, sign_data, aclr,
                        result, cout, overflow);
    parameter width_in = 4;     
    parameter width_out = 8;    
    parameter lpm_representation = "UNSIGNED";
    parameter extra_latency = 0;
    parameter use_wys = "ON";
    parameter lpm_hint = "UNUSED";
    parameter lpm_type = "altaccumulate";
    input cin;
    input [width_in-1:0] data;  
    input add_sub;              
    input clock;                
    input sload;                
    input clken;                
    input sign_data;            
    input aclr;                 
    output [width_out-1:0] result;  
    output cout;
    output overflow;
    reg [width_out:0] temp_sum;
    reg overflow;
    reg overflow_int;
    reg cout_int;
    reg cout_delayed;
    reg [width_out-1:0] result;
    reg [width_out+1:0] result_int;
    reg [(width_out - width_in) : 0] zeropad;
    reg borrow;
    reg cin_int;
    reg [width_out-1:0] fb_int;
    reg [width_out -1:0] data_int;
    reg [width_out+1:0] result_pipe [extra_latency:0];
    reg [width_out+1:0] result_full;
    reg [width_out+1:0] result_full2;
    reg a;
    wire [width_out:0] temp_sum_wire;
    wire cout;
    wire cout_int_wire;
    wire cout_delayed_wire;
    wire overflow_int_wire;
    wire [width_out+1:0] result_int_wire;
    tri0 aclr_int;
    tri0 sign_data_int;
    tri0 sload_int;
    tri1 clken_int;
    tri1 add_sub_int;
    integer head;
    integer i;
    initial
    begin
        if( width_in <= 0 )
        begin
            $display("Error! Value of width_in parameter must be greater than 0.");
            $stop;
        end
        if( width_out <= 0 )
        begin
            $display("Error! Value of width_out parameter must be greater than 0.");
            $stop;
        end
        if( extra_latency > width_out )
        begin
            $display("Info: Value of extra_latency parameter should be lower than width_out parameter for better performance/utilization.");
        end
        if( width_in > width_out )
        begin
            $display("Error! Value of width_in parameter should be lower than or equal to width_out.");
            $stop;
        end
        result = 0;
        cout_delayed = 0;
        overflow = 0;
        head = 0;
        result_int = 0;
        for (i = 0; i <= extra_latency; i = i +1)
        begin
            result_pipe [i] = 0;
        end
    end
    always @(posedge clock or posedge aclr_int)
    begin
        if (aclr_int == 1)
        begin
            result_int = 0;
            result = 0;
            overflow = 0;
            cout_delayed = 0;
            for (i = 0; i <= extra_latency; i = i +1)
            begin
                result_pipe [i] = 0;
            end
        end
        else
        begin
            if (clken_int == 1)
            begin
                if (extra_latency > 0)
                begin
                    result_pipe [head] = {
                                            result_int [width_out+1],
                                            {cout_int_wire, result_int [width_out-1:0]}
                                        };
                    head = (head + 1) % (extra_latency);
                    result_full = result_pipe [head];
                    cout_delayed = result_full [width_out];
                    result = result_full [width_out-1:0];
                    overflow = result_full [width_out+1];
                end
                else
                begin
                    result = temp_sum_wire;
                    overflow = overflow_int_wire;
                end
                result_int = {overflow_int_wire, {cout_int_wire, temp_sum_wire [width_out-1:0]}};
            end
        end
    end
    always @ (data or cin or add_sub_int or sign_data_int or
                result_int_wire [width_out -1:0] or sload_int)
    begin
        if ((lpm_representation == "SIGNED") || (sign_data_int == 1))
        begin
            zeropad = (data [width_in-1] ==0) ? 0 : -1;
        end
        else
        begin
            zeropad = 0;
        end
        fb_int = (sload_int == 1'b1) ? 0 : result_int_wire [width_out-1:0];
        data_int = {zeropad, data};
        if ((add_sub_int == 1) || (sload_int == 1))
        begin
            cin_int = ((sload_int == 1'b1) ? 0 : ((cin === 1'bz) ? 0 : cin));
            temp_sum = fb_int + data_int + cin_int;
            cout_int = temp_sum [width_out];
        end
        else
        begin
            cin_int = (cin === 1'bz) ? 1 : cin;
            borrow = ~cin_int;
            temp_sum = fb_int - data_int - borrow;
            result_full2 = data_int + borrow;
            cout_int = (fb_int >= result_full2) ? 1 : 0;
        end
        if ((lpm_representation == "SIGNED") || (sign_data_int == 1))
        begin
            a = (data [width_in-1] ~^ fb_int [width_out-1]) ^ (~add_sub_int);
            overflow_int = a & (fb_int [width_out-1] ^ temp_sum[width_out-1]);
        end
        else
        begin
            overflow_int = (add_sub_int == 1) ? cout_int : ~cout_int;
        end
        if (sload_int == 1)
        begin
            cout_int = !add_sub_int;
            overflow_int = 0;
        end
    end
    assign sign_data_int = sign_data;
    assign sload_int =  sload;
    assign add_sub_int = add_sub;
    assign clken_int = clken;
    assign aclr_int = aclr;
    assign result_int_wire = result_int;
    assign temp_sum_wire = temp_sum;
    assign cout_int_wire = cout_int;
    assign overflow_int_wire = overflow_int;
    assign cout = (extra_latency == 0) ? cout_int_wire : cout_delayed_wire;
    assign cout_delayed_wire = cout_delayed;
endmodule




 `timescale 1ns / 1ps

module tb;

    // Parameters
    parameter WIDTH_IN = 4;
    parameter WIDTH_OUT = 8;

    // Testbench signals
    reg cin;
    reg [WIDTH_IN-1:0] data;
    reg add_sub;
    reg clock;
    reg sload;
    reg clken;
    reg sign_data;
    reg aclr;
    
    // Outputs
    wire [WIDTH_OUT-1:0] result_ref, result_dut;
    wire cout_ref, cout_dut;
    wire overflow_ref, overflow_dut;

    wire match;

    integer total_tests = 0;
	integer failed_tests = 0;

    assign match = ({result_ref, cout_ref, overflow_ref} === ({result_ref, cout_ref, overflow_ref} ^ {result_dut, cout_dut, overflow_dut} ^ {result_ref, cout_ref, overflow_ref}));


    // Instantiate the altaccumulate module
    altaccumulate_ref #(
        .width_in(WIDTH_IN),
        .width_out(WIDTH_OUT),
        .extra_latency(1)
    ) ref_model (
        .cin(cin),
        .data(data),
        .add_sub(add_sub),
        .clock(clock),
        .sload(sload),
        .clken(clken),
        .sign_data(sign_data),
        .aclr(aclr),
        .result(result_ref),
        .cout(cout_ref),
        .overflow(overflow_ref)
    );

    altaccumulate #(
        .width_in(WIDTH_IN),
        .width_out(WIDTH_OUT),
        .extra_latency(1)
    ) uut (
        .cin(cin),
        .data(data),
        .add_sub(add_sub),
        .clock(clock),
        .sload(sload),
        .clken(clken),
        .sign_data(sign_data),
        .aclr(aclr),
        .result(result_dut),
        .cout(cout_dut),
        .overflow(overflow_dut)
    );


    // Clock generation
    initial begin
        clock = 0;
        forever #5 clock = ~clock; // 100 MHz clock
    end

    // Test procedure
    initial begin
        // Initialize signals
        cin = 0;
        data = 0;
        add_sub = 0;
        sload = 0;
        clken = 0;
        sign_data = 0;
        aclr = 0;

        // Release reset
        #10;
        aclr = 1; // Assert reset
        #10;
        aclr = 0;// De-assert reset
        clken = 1;

        //Load
        @(negedge clock);
        sload = 1;
        data = 4'hA;
        @(negedge clock);
        sign_data = 1;
        add_sub = 0;
        sload = 0;
        data = 4'hF;
        cin = 0;
        @(negedge clock);
        compare();

        
        // Test Case 1: Addition
        repeat (25) begin
            data = $random; // Input data
            add_sub = 1; // Addition
            cin = $random; // Carry in
            sload = 0; // Not loading
            @(negedge clock);
            compare();
        end

        @(negedge clock);
        compare();
        sload = 1;
        data = 4'hF;
        @(negedge clock);
        compare();

        // Test Case 2: Subtraction
        repeat (25) begin
            data = $random; // Input data
            add_sub = 0; // Addition
            cin = $random; // Carry in
            sload = 0; // Not loading
            @(negedge clock);
            compare();
        end

        @(negedge clock);
        compare();
        sload = 1;
        data = 4'h7;
        @(negedge clock);
        compare();
        sload = 0; // Not loading

        
        repeat (45) begin
            data = $random; // Input data
            add_sub = $random; // Addition
            cin = $random; // Carry in
            sign_data = $random;
            @(negedge clock);
            compare();
        end

        #10;
        aclr = 1; // Assert reset
        clken = 0;
        #10;
        aclr = 0;// De-assert reset
        clken = 1;
        $display("\033[1;34mTotal testcases: %d, Failed testcases: %d\033[0m", total_tests, failed_tests);
        if (failed_tests==0) begin
            $display("=====================Your Design Passed======================");
    end
        // Finish simulation
        $finish;
    end

    task compare;
    begin
        total_tests = total_tests + 1;

        if (match)                                //condition to check DUT outputs and calculated 
                                                    //outputs from task are equal 
			begin
			//	$display("\033[1;32mtestcase is passed!!!\033[0m");
//				$display("testcase is passed!!!");
           // 	$display("cin, data = %h, add_sub = %h, sload = %h, clken = %h, sign_data = %h, aclr = %h, result_dut = %h, cout_dut = %h, overflow_dut = %h, result_ref = %h, cout_ref = %h, overflow_ref = %h", cin, data, add_sub, sload, clken, sign_data, aclr, result_dut, cout_dut, overflow_dut, result_ref, cout_ref, overflow_ref);      //displaying inputs, outputs and result
			end

		else begin
		//	$display("\033[1;31mtestcase is failed!!!\033[0m");
         //   $display("cin, data = %h, add_sub = %h, sload = %h, clken = %h, sign_data = %h, aclr = %h, result_dut = %h, cout_dut = %h, overflow_dut = %h, result_ref = %h, cout_ref = %h, overflow_ref = %h", cin, data, add_sub, sload, clken, sign_data, aclr, result_dut, cout_dut, overflow_dut, result_ref, cout_ref, overflow_ref);      //displaying inputs, outputs and result
            failed_tests = failed_tests + 1; 
		end
    end
	endtask


    initial begin
        $dumpfile("sim.fsdb");
        $dumpvars(0);
    end
    
endmodule
