 
module ref_eth_cop
(
  wb_clk_i, wb_rst_i, 
  m1_wb_adr_i, m1_wb_sel_i, m1_wb_we_i,  ref_m1_wb_dat_o, 
  m1_wb_dat_i, m1_wb_cyc_i, m1_wb_stb_i, ref_m1_wb_ack_o, 
  ref_m1_wb_err_o, 
  m2_wb_adr_i, m2_wb_sel_i, m2_wb_we_i,  ref_m2_wb_dat_o, 
  m2_wb_dat_i, m2_wb_cyc_i, m2_wb_stb_i, ref_m2_wb_ack_o, 
  ref_m2_wb_err_o, 
 	ref_s1_wb_adr_o, ref_s1_wb_sel_o, ref_s1_wb_we_o,  ref_s1_wb_cyc_o, 
 	ref_s1_wb_stb_o, s1_wb_ack_i, s1_wb_err_i, s1_wb_dat_i,
 	ref_s1_wb_dat_o, 
 	ref_s2_wb_adr_o, ref_s2_wb_sel_o, ref_s2_wb_we_o,  ref_s2_wb_cyc_o, 
 	ref_s2_wb_stb_o, s2_wb_ack_i, s2_wb_err_i, s2_wb_dat_i,
 	ref_s2_wb_dat_o
);
parameter ETH_BASE     = 32'hd0000000;
parameter ETH_WIDTH    = 32'h800;
parameter MEMORY_BASE  = 32'h2000;
parameter MEMORY_WIDTH = 32'h10000;
input wb_clk_i, wb_rst_i;
input  [31:0] m1_wb_adr_i, m1_wb_dat_i;
input   [3:0] m1_wb_sel_i;
input         m1_wb_cyc_i, m1_wb_stb_i, m1_wb_we_i;
output [31:0] ref_m1_wb_dat_o;
output        ref_m1_wb_ack_o, ref_m1_wb_err_o;
input  [31:0] m2_wb_adr_i, m2_wb_dat_i;
input   [3:0] m2_wb_sel_i;
input         m2_wb_cyc_i, m2_wb_stb_i, m2_wb_we_i;
output [31:0] ref_m2_wb_dat_o;
output        ref_m2_wb_ack_o, ref_m2_wb_err_o;
input  [31:0] s1_wb_dat_i;
input         s1_wb_ack_i, s1_wb_err_i;
output [31:0] ref_s1_wb_adr_o, ref_s1_wb_dat_o;
output  [3:0] ref_s1_wb_sel_o;
output        ref_s1_wb_we_o,  ref_s1_wb_cyc_o, ref_s1_wb_stb_o;
input  [31:0] s2_wb_dat_i;
input         s2_wb_ack_i, s2_wb_err_i;
output [31:0] ref_s2_wb_adr_o, ref_s2_wb_dat_o;
output  [3:0] ref_s2_wb_sel_o;
output        ref_s2_wb_we_o,  ref_s2_wb_cyc_o, ref_s2_wb_stb_o;
reg           m1_in_progress;
reg           m2_in_progress;
reg    [31:0] ref_s1_wb_adr_o;
reg     [3:0] ref_s1_wb_sel_o;
reg           ref_s1_wb_we_o;
reg    [31:0] ref_s1_wb_dat_o;
reg           ref_s1_wb_cyc_o;
reg           ref_s1_wb_stb_o;
reg    [31:0] ref_s2_wb_adr_o;
reg     [3:0] ref_s2_wb_sel_o;
reg           ref_s2_wb_we_o;
reg    [31:0] ref_s2_wb_dat_o;
reg           ref_s2_wb_cyc_o;
reg           ref_s2_wb_stb_o;
reg           ref_m1_wb_ack_o;
reg    [31:0] ref_m1_wb_dat_o;
reg           ref_m2_wb_ack_o;
reg    [31:0] ref_m2_wb_dat_o;
reg           ref_m1_wb_err_o;
reg           ref_m2_wb_err_o;
wire m_wb_access_finished;
wire m1_addressed_s1 = (m1_wb_adr_i >= ETH_BASE) &
                       (m1_wb_adr_i < (ETH_BASE + ETH_WIDTH));
wire m1_addressed_s2 = (m1_wb_adr_i >= MEMORY_BASE) &
                       (m1_wb_adr_i < (MEMORY_BASE + MEMORY_WIDTH));
wire m2_addressed_s1 = (m2_wb_adr_i >= ETH_BASE) &
                       (m2_wb_adr_i < (ETH_BASE + ETH_WIDTH));
wire m2_addressed_s2 = (m2_wb_adr_i >= MEMORY_BASE) &
                       (m2_wb_adr_i < (MEMORY_BASE + MEMORY_WIDTH));
wire m1_req = m1_wb_cyc_i & m1_wb_stb_i & (m1_addressed_s1 | m1_addressed_s2);
wire m2_req = m2_wb_cyc_i & m2_wb_stb_i & (m2_addressed_s1 | m2_addressed_s2);
always @ (posedge wb_clk_i or posedge wb_rst_i)
begin
  if(wb_rst_i)
    begin
      m1_in_progress <= 0;
      m2_in_progress <= 0;
      ref_s1_wb_adr_o    <= 0;
      ref_s1_wb_sel_o    <= 0;
      ref_s1_wb_we_o     <= 0;
      ref_s1_wb_dat_o    <= 0;
      ref_s1_wb_cyc_o    <= 0;
      ref_s1_wb_stb_o    <= 0;
      ref_s2_wb_adr_o    <= 0;
      ref_s2_wb_sel_o    <= 0;
      ref_s2_wb_we_o     <= 0;
      ref_s2_wb_dat_o    <= 0;
      ref_s2_wb_cyc_o    <= 0;
      ref_s2_wb_stb_o    <= 0;
    end
  else
    begin
      case({m1_in_progress, m2_in_progress, m1_req, m2_req, m_wb_access_finished})  
        5'b00_10_0, 5'b00_11_0 :
          begin
            m1_in_progress <= 1'b1;  
            if(m1_addressed_s1)
              begin
                ref_s1_wb_adr_o <= m1_wb_adr_i;
                ref_s1_wb_sel_o <= m1_wb_sel_i;
                ref_s1_wb_we_o  <= m1_wb_we_i;
                ref_s1_wb_dat_o <= m1_wb_dat_i;
                ref_s1_wb_cyc_o <= 1'b1;
                ref_s1_wb_stb_o <= 1'b1;
              end
            else if(m1_addressed_s2)
              begin
                ref_s2_wb_adr_o <= m1_wb_adr_i;
                ref_s2_wb_sel_o <= m1_wb_sel_i;
                ref_s2_wb_we_o  <= m1_wb_we_i;
                ref_s2_wb_dat_o <= m1_wb_dat_i;
                ref_s2_wb_cyc_o <= 1'b1;
                ref_s2_wb_stb_o <= 1'b1;
              end
            else
              $display("(%t)(%m)WISHBONE ERROR: Unspecified address space accessed", $time);
          end
        5'b00_01_0 :
          begin
            m2_in_progress <= 1'b1;  
            if(m2_addressed_s1)
              begin
                ref_s1_wb_adr_o <= m2_wb_adr_i;
                ref_s1_wb_sel_o <= m2_wb_sel_i;
                ref_s1_wb_we_o  <= m2_wb_we_i;
                ref_s1_wb_dat_o <= m2_wb_dat_i;
                ref_s1_wb_cyc_o <= 1'b1;
                ref_s1_wb_stb_o <= 1'b1;
              end
            else if(m2_addressed_s2)
              begin
                ref_s2_wb_adr_o <= m2_wb_adr_i;
                ref_s2_wb_sel_o <= m2_wb_sel_i;
                ref_s2_wb_we_o  <= m2_wb_we_i;
                ref_s2_wb_dat_o <= m2_wb_dat_i;
                ref_s2_wb_cyc_o <= 1'b1;
                ref_s2_wb_stb_o <= 1'b1;
              end
            else
              $display("(%t)(%m)WISHBONE ERROR: Unspecified address space accessed", $time);
          end
        5'b10_10_1, 5'b10_11_1 :
          begin
            m1_in_progress <= 1'b0;  
            if(m1_addressed_s1)
              begin
                ref_s1_wb_cyc_o <= 1'b0;
                ref_s1_wb_stb_o <= 1'b0;
              end
            else if(m1_addressed_s2)
              begin
                ref_s2_wb_cyc_o <= 1'b0;
                ref_s2_wb_stb_o <= 1'b0;
              end
          end
        5'b01_01_1, 5'b01_11_1 :
          begin
            m2_in_progress <= 1'b0;  
            if(m2_addressed_s1)
              begin
                ref_s1_wb_cyc_o <= 1'b0;
                ref_s1_wb_stb_o <= 1'b0;
              end
            else if(m2_addressed_s2)
              begin
                ref_s2_wb_cyc_o <= 1'b0;
                ref_s2_wb_stb_o <= 1'b0;
              end
          end
      endcase
    end
end
always @ (m1_in_progress or m1_wb_adr_i or s1_wb_ack_i or s2_wb_ack_i or s1_wb_dat_i or s2_wb_dat_i or m1_addressed_s1 or m1_addressed_s2)
begin
  if(m1_in_progress)
    begin
      if(m1_addressed_s1) begin
        ref_m1_wb_ack_o <= s1_wb_ack_i;
        ref_m1_wb_dat_o <= s1_wb_dat_i;
      end
      else if(m1_addressed_s2) begin
        ref_m1_wb_ack_o <= s2_wb_ack_i;
        ref_m1_wb_dat_o <= s2_wb_dat_i;
      end
    end
  else
    ref_m1_wb_ack_o <= 0;
end
always @ (m2_in_progress or m2_wb_adr_i or s1_wb_ack_i or s2_wb_ack_i or s1_wb_dat_i or s2_wb_dat_i or m2_addressed_s1 or m2_addressed_s2)
begin
  if(m2_in_progress)
    begin
      if(m2_addressed_s1) begin
        ref_m2_wb_ack_o <= s1_wb_ack_i;
        ref_m2_wb_dat_o <= s1_wb_dat_i;
      end
      else if(m2_addressed_s2) begin
        ref_m2_wb_ack_o <= s2_wb_ack_i;
        ref_m2_wb_dat_o <= s2_wb_dat_i;
      end
    end
  else
    ref_m2_wb_ack_o <= 0;
end
always @ (m1_in_progress or m1_wb_adr_i or s1_wb_err_i or s2_wb_err_i or m2_addressed_s1 or m2_addressed_s2 or
          m1_wb_cyc_i or m1_wb_stb_i)
begin
  if(m1_in_progress)  begin
    if(m1_addressed_s1)
      ref_m1_wb_err_o <= s1_wb_err_i;
    else if(m1_addressed_s2)
      ref_m1_wb_err_o <= s2_wb_err_i;
  end
  else if(m1_wb_cyc_i & m1_wb_stb_i & ~m1_addressed_s1 & ~m1_addressed_s2)
    ref_m1_wb_err_o <= 1'b1;
  else
    ref_m1_wb_err_o <= 1'b0;
end
always @ (m2_in_progress or m2_wb_adr_i or s1_wb_err_i or s2_wb_err_i or m2_addressed_s1 or m2_addressed_s2 or
          m2_wb_cyc_i or m2_wb_stb_i)
begin
  if(m2_in_progress)  begin
    if(m2_addressed_s1)
      ref_m2_wb_err_o <= s1_wb_err_i;
    else if(m2_addressed_s2)
      ref_m2_wb_err_o <= s2_wb_err_i;
  end
  else if(m2_wb_cyc_i & m2_wb_stb_i & ~m2_addressed_s1 & ~m2_addressed_s2)
    ref_m2_wb_err_o <= 1'b1;
  else
    ref_m2_wb_err_o <= 1'b0;
end
assign m_wb_access_finished = ref_m1_wb_ack_o | ref_m1_wb_err_o | ref_m2_wb_ack_o | ref_m2_wb_err_o;
integer cnt;
always @ (posedge wb_clk_i or posedge wb_rst_i)
begin
  if(wb_rst_i)
    cnt <= 0;
  else
  if(s1_wb_ack_i | s1_wb_err_i | s2_wb_ack_i | s2_wb_err_i)
    cnt <= 0;
  else
  if(ref_s1_wb_cyc_o | ref_s2_wb_cyc_o)
    cnt <= cnt+1;
end
always @ (posedge wb_clk_i)
begin
  if(cnt==1000) begin
    $display("(%0t)(%m) ERROR: WB activity ??? ", $time);
    if(ref_s1_wb_cyc_o) begin
      $display("ref_s1_wb_dat_o = 0x%0x", ref_s1_wb_dat_o);
      $display("ref_s1_wb_adr_o = 0x%0x", ref_s1_wb_adr_o);
      $display("ref_s1_wb_sel_o = 0x%0x", ref_s1_wb_sel_o);
      $display("ref_s1_wb_we_o = 0x%0x", ref_s1_wb_we_o);
    end
    else if(ref_s2_wb_cyc_o) begin
      $display("ref_s2_wb_dat_o = 0x%0x", ref_s2_wb_dat_o);
      $display("ref_s2_wb_adr_o = 0x%0x", ref_s2_wb_adr_o);
      $display("ref_s2_wb_sel_o = 0x%0x", ref_s2_wb_sel_o);
      $display("ref_s2_wb_we_o = 0x%0x", ref_s2_wb_we_o);
    end
    $stop;
  end
end
always @ (posedge wb_clk_i)
begin
  if(s1_wb_err_i & ref_s1_wb_cyc_o) begin
    $display("(%0t) ERROR: WB cycle finished with error acknowledge ", $time);
    $display("ref_s1_wb_dat_o = 0x%0x", ref_s1_wb_dat_o);
    $display("ref_s1_wb_adr_o = 0x%0x", ref_s1_wb_adr_o);
    $display("ref_s1_wb_sel_o = 0x%0x", ref_s1_wb_sel_o);
    $display("ref_s1_wb_we_o = 0x%0x", ref_s1_wb_we_o);
    $stop;
  end
  if(s2_wb_err_i & ref_s2_wb_cyc_o) begin
    $display("(%0t) ERROR: WB cycle finished with error acknowledge ", $time);
    $display("ref_s2_wb_dat_o = 0x%0x", ref_s2_wb_dat_o);
    $display("ref_s2_wb_adr_o = 0x%0x", ref_s2_wb_adr_o);
    $display("ref_s2_wb_sel_o = 0x%0x", ref_s2_wb_sel_o);
    $display("ref_s2_wb_we_o = 0x%0x", ref_s2_wb_we_o);
    $stop;
  end
end
endmodule




 `timescale 1ns / 1ps

module tb;

    // Parameters
    parameter CLK_PERIOD = 10; // Clock period for wb_clk_i

    // Inputs
    reg wb_clk_i;
    reg wb_rst_i;
    reg [31:0] m1_wb_adr_i, m1_wb_dat_i;
    reg [3:0] m1_wb_sel_i;
    reg m1_wb_cyc_i, m1_wb_stb_i, m1_wb_we_i;
    reg [31:0] m2_wb_adr_i, m2_wb_dat_i;
    reg [3:0] m2_wb_sel_i;
    reg m2_wb_cyc_i, m2_wb_stb_i, m2_wb_we_i;
    reg [31:0] s1_wb_dat_i, s2_wb_dat_i;
    reg s1_wb_ack_i, s1_wb_err_i;
    reg s2_wb_ack_i, s2_wb_err_i;

    // ref Outputs
    wire [31:0] ref_m1_wb_dat_o;
    wire ref_m1_wb_ack_o, ref_m1_wb_err_o;
    wire [31:0] ref_m2_wb_dat_o;
    wire ref_m2_wb_ack_o, ref_m2_wb_err_o;
    wire [31:0] ref_s1_wb_adr_o, ref_s1_wb_dat_o;
    wire [3:0] ref_s1_wb_sel_o;
    wire ref_s1_wb_we_o, ref_s1_wb_cyc_o, ref_s1_wb_stb_o;
    wire [31:0] ref_s2_wb_adr_o, ref_s2_wb_dat_o;
    wire [3:0] ref_s2_wb_sel_o;
    wire ref_s2_wb_we_o, ref_s2_wb_cyc_o, ref_s2_wb_stb_o;

    // Outputs
    wire [31:0] m1_wb_dat_o;
    wire m1_wb_ack_o, m1_wb_err_o;
    wire [31:0] m2_wb_dat_o;
    wire m2_wb_ack_o, m2_wb_err_o;
    wire [31:0] s1_wb_adr_o, s1_wb_dat_o;
    wire [3:0] s1_wb_sel_o;
    wire s1_wb_we_o, s1_wb_cyc_o, s1_wb_stb_o;
    wire [31:0] s2_wb_adr_o, s2_wb_dat_o;
    wire [3:0] s2_wb_sel_o;
    wire s2_wb_we_o, s2_wb_cyc_o, s2_wb_stb_o;

	wire match;
 	integer total_tests = 0;
	integer failed_tests = 0;

assign match = ({ref_m1_wb_dat_o,ref_m1_wb_ack_o, ref_m1_wb_err_o,ref_m2_wb_dat_o,ref_m2_wb_ack_o, ref_m2_wb_err_o,ref_s1_wb_adr_o, ref_s1_wb_dat_o,ref_s1_wb_sel_o,ref_s1_wb_we_o, ref_s1_wb_cyc_o, ref_s1_wb_stb_o,ref_s2_wb_adr_o, ref_s2_wb_dat_o,ref_s2_wb_sel_o,ref_s2_wb_we_o, ref_s2_wb_cyc_o, ref_s2_wb_stb_o} === {m1_wb_dat_o,m1_wb_ack_o, m1_wb_err_o,m2_wb_dat_o,m2_wb_ack_o, m2_wb_err_o,s1_wb_adr_o,s1_wb_dat_o,s1_wb_sel_o,s1_wb_we_o, s1_wb_cyc_o, s1_wb_stb_o,s2_wb_adr_o, s2_wb_dat_o,s2_wb_sel_o,s2_wb_we_o,ref_s2_wb_cyc_o, s2_wb_stb_o} );

    // Instantiate the eth_cop module
    ref_eth_cop rf(
        .wb_clk_i(wb_clk_i),
        .wb_rst_i(wb_rst_i),
        .m1_wb_adr_i(m1_wb_adr_i), .m1_wb_dat_i(m1_wb_dat_i),
        .m1_wb_sel_i(m1_wb_sel_i), .m1_wb_cyc_i(m1_wb_cyc_i),
        .m1_wb_stb_i(m1_wb_stb_i), .m1_wb_we_i(m1_wb_we_i),
        .ref_m1_wb_dat_o(ref_m1_wb_dat_o), .ref_m1_wb_ack_o(ref_m1_wb_ack_o),
        .ref_m1_wb_err_o(ref_m1_wb_err_o),
        .m2_wb_adr_i(m2_wb_adr_i), .m2_wb_dat_i(m2_wb_dat_i),
        .m2_wb_sel_i(m2_wb_sel_i), .m2_wb_cyc_i(m2_wb_cyc_i),
        .m2_wb_stb_i(m2_wb_stb_i), .m2_wb_we_i(m2_wb_we_i),
        .ref_m2_wb_dat_o(ref_m2_wb_dat_o), .ref_m2_wb_ack_o(ref_m2_wb_ack_o),
        .ref_m2_wb_err_o(ref_m2_wb_err_o),
        .ref_s1_wb_adr_o(ref_s1_wb_adr_o), .ref_s1_wb_dat_o(ref_s1_wb_dat_o),
        .ref_s1_wb_sel_o(ref_s1_wb_sel_o), .ref_s1_wb_we_o(ref_s1_wb_we_o),
        .ref_s1_wb_cyc_o(ref_s1_wb_cyc_o), .ref_s1_wb_stb_o(ref_s1_wb_stb_o),
        .s1_wb_ack_i(s1_wb_ack_i), .s1_wb_err_i(s1_wb_err_i),
        .s1_wb_dat_i(s1_wb_dat_i),
        .ref_s2_wb_adr_o(ref_s2_wb_adr_o), .ref_s2_wb_dat_o(ref_s2_wb_dat_o),
        .ref_s2_wb_sel_o(ref_s2_wb_sel_o), .ref_s2_wb_we_o(ref_s2_wb_we_o),
        .ref_s2_wb_cyc_o(ref_s2_wb_cyc_o), .ref_s2_wb_stb_o(ref_s2_wb_stb_o),
        .s2_wb_ack_i(s2_wb_ack_i), .s2_wb_err_i(s2_wb_err_i),
        .s2_wb_dat_i(s2_wb_dat_i)
    );

    // Instantiate the eth_cop module
   eth_cop dut (
        .wb_clk_i(wb_clk_i),
        .wb_rst_i(wb_rst_i),
        .m1_wb_adr_i(m1_wb_adr_i), .m1_wb_dat_i(m1_wb_dat_i),
        .m1_wb_sel_i(m1_wb_sel_i), .m1_wb_cyc_i(m1_wb_cyc_i),
        .m1_wb_stb_i(m1_wb_stb_i), .m1_wb_we_i(m1_wb_we_i),
        .m1_wb_dat_o(m1_wb_dat_o), .m1_wb_ack_o(m1_wb_ack_o),
        .m1_wb_err_o(m1_wb_err_o),
        .m2_wb_adr_i(m2_wb_adr_i), .m2_wb_dat_i(m2_wb_dat_i),
        .m2_wb_sel_i(m2_wb_sel_i), .m2_wb_cyc_i(m2_wb_cyc_i),
        .m2_wb_stb_i(m2_wb_stb_i), .m2_wb_we_i(m2_wb_we_i),
        .m2_wb_dat_o(m2_wb_dat_o), .m2_wb_ack_o(m2_wb_ack_o),
        .m2_wb_err_o(m2_wb_err_o),
        .s1_wb_adr_o(s1_wb_adr_o), .s1_wb_dat_o(s1_wb_dat_o),
        .s1_wb_sel_o(s1_wb_sel_o), .s1_wb_we_o(s1_wb_we_o),
        .s1_wb_cyc_o(s1_wb_cyc_o), .s1_wb_stb_o(s1_wb_stb_o),
        .s1_wb_ack_i(s1_wb_ack_i), .s1_wb_err_i(s1_wb_err_i),
        .s1_wb_dat_i(s1_wb_dat_i),
        .s2_wb_adr_o(s2_wb_adr_o), .s2_wb_dat_o(s2_wb_dat_o),
        .s2_wb_sel_o(s2_wb_sel_o), .s2_wb_we_o(s2_wb_we_o),
        .s2_wb_cyc_o(s2_wb_cyc_o), .s2_wb_stb_o(s2_wb_stb_o),
        .s2_wb_ack_i(s2_wb_ack_i), .s2_wb_err_i(s2_wb_err_i),
        .s2_wb_dat_i(s2_wb_dat_i)
    );

    // Generate clock signal
    initial begin
        wb_clk_i = 0;
        forever #(CLK_PERIOD / 2) wb_clk_i = ~wb_clk_i; // Toggle clock
    end

    // Test Procedure
    initial begin
        // Initialize inputs
        wb_rst_i = 1;
        m1_wb_adr_i = 0; m1_wb_dat_i = 0; m1_wb_sel_i = 0;
        m1_wb_cyc_i = 0; m1_wb_stb_i = 0; m1_wb_we_i = 0;
        m2_wb_adr_i = 0; m2_wb_dat_i = 0; m2_wb_sel_i = 0;
        m2_wb_cyc_i = 0; m2_wb_stb_i = 0; m2_wb_we_i = 0;
        s1_wb_dat_i = 0; s2_wb_dat_i = 0;
        s1_wb_ack_i = 0; s1_wb_err_i = 0;
        s2_wb_ack_i = 0; s2_wb_err_i = 0;

        // Apply reset
        #(CLK_PERIOD);
        wb_rst_i = 0; // De-assert reset
        #(CLK_PERIOD);

        // Test Case 1: Simple Write to s1
        m1_wb_adr_i = 32'hd0000000; // Address for s1
        m1_wb_dat_i = 32'hA5A5A5A5; // Data to write
        m1_wb_sel_i = 4'b1111; // Select all bytes
        m1_wb_cyc_i = 1; // Assert cycle
        m1_wb_stb_i = 1; // Assert strobe
        m1_wb_we_i = 1; // Write enable
        #(CLK_PERIOD);
        m1_wb_cyc_i = 0; // End cycle
        m1_wb_stb_i = 0; // End strobe
        #(CLK_PERIOD);
compare();

        // Test Case 2: Read from s1
        s1_wb_ack_i = 1; // Simulate acknowledgment from slave
        s1_wb_dat_i = 32'hA5A5A5A5; // Simulated data from slave
        m1_wb_adr_i = 32'hd0000000; // Address for s1
        m1_wb_cyc_i = 1; // Assert cycle
        m1_wb_stb_i = 1; // Assert strobe
        m1_wb_we_i = 0; // Read
        #(CLK_PERIOD);
        m1_wb_cyc_i = 0; // End cycle
        m1_wb_stb_i = 0; // End strobe
        #(CLK_PERIOD);
compare();

        // Test Case 3: Write to s2
        m2_wb_adr_i = 32'h2000; // Address for s2
        m2_wb_dat_i = 32'h5A5A5A5A; // Data to write
        m2_wb_sel_i = 4'b1111; // Select all bytes
        m2_wb_cyc_i = 1; // Assert cycle
        m2_wb_stb_i = 1; // Assert strobe
        m2_wb_we_i = 1; // Write enable
        #(CLK_PERIOD);
        m2_wb_cyc_i = 0; // End cycle
        m2_wb_stb_i = 0; // End strobe
        #(CLK_PERIOD);

compare();

        // Test Case 4: Read from s2
        s2_wb_ack_i = 1; // Simulate acknowledgment from slave
        s2_wb_dat_i = 32'h5A5A5A5A; // Simulated data from slave
        m2_wb_adr_i = 32'h2000; // Address for s2
        m2_wb_cyc_i = 1; // Assert cycle
        m2_wb_stb_i = 1; // Assert strobe
        m2_wb_we_i = 0; // Read
        #(CLK_PERIOD);
        m2_wb_cyc_i = 0; // End cycle
        m2_wb_stb_i = 0; // End strobe
        #(CLK_PERIOD);
compare();
 

repeat (1000) begin
            @(negedge wb_clk_i);
	m1_wb_adr_i = $random;
	m1_wb_dat_i = $random;
	m1_wb_sel_i = $random;
	m1_wb_cyc_i = $random;
	m1_wb_stb_i = $random;
	m1_wb_we_i = $random;
	m2_wb_adr_i = $random;
	m2_wb_dat_i = $random;
	m2_wb_sel_i = $random;
	m2_wb_cyc_i = $random;
	m2_wb_stb_i = $random;
	m2_wb_we_i = $random;
	s1_wb_dat_i = $random;
	s2_wb_dat_i = $random;
	s1_wb_ack_i = $random;
	s1_wb_err_i = $random;
	s2_wb_ack_i = $random;
	s2_wb_err_i = $random;
compare();
end
 	$display("All tests passed: design passed");
        $display("\033[1;34mTotal testcases: %d, Failed testcases: %d\033[0m", total_tests, failed_tests);
        // Finish simulation

    if (failed_tests==0) begin
            $display("=====================Your Design Passed======================");
    end
        #(CLK_PERIOD * 10);
        $finish;
    end

task compare;
        total_tests = total_tests + 1;
        if (match)                                //condition to check DUT outputs and calculated 
                                                    //outputs from task are equal 
			begin
				//$display("\033[1;32mtestcase is passed!!!\033[0m");
			end

		else begin
			//$display("\033[1;31mtestcase is failed!!!\033[0m");
            failed_tests = failed_tests + 1; 
		end
    
	endtask
endmodule
