 

module ref_aeMB_xecu (
   ref_dwb_adr_o, ref_dwb_sel_o, ref_fsl_adr_o, ref_fsl_tag_o, ref_rRESULT, ref_rDWBSEL,
   ref_rMSR_IE, ref_rMSR_BIP,
   rREGA, rREGB, rMXSRC, rMXTGT, rRA, rRB, rMXALU, rBRA, rDLY, rALT,
   rSTALL, rSIMM, rIMM, rOPC, rRD, rDWBDI, rPC, gclk, grst, gena
   );
   parameter DW=32;
   parameter MUL=0;
   parameter BSF=0;   
   output [DW-1:2] ref_dwb_adr_o;
   output [3:0]    ref_dwb_sel_o;
   output [6:2]   ref_fsl_adr_o;
   output [1:0]   ref_fsl_tag_o;   
   output [31:0]   ref_rRESULT;
   output [3:0]    ref_rDWBSEL;   
   output 	   ref_rMSR_IE;
   output 	   ref_rMSR_BIP;
   input [31:0]    rREGA, rREGB;
   input [1:0] 	   rMXSRC, rMXTGT;
   input [4:0] 	   rRA, rRB;
   input [2:0] 	   rMXALU;
   input 	   rBRA, rDLY;
   input [10:0]    rALT;   
   input 	   rSTALL;   
   input [31:0]    rSIMM;
   input [15:0]    rIMM;
   input [5:0] 	   rOPC;
   input [4:0] 	   rRD;   
   input [31:0]    rDWBDI;
   input [31:2]    rPC;   
   input 	   gclk, grst, gena;
   reg 		   rMSR_C, xMSR_C;
   reg 		   ref_rMSR_IE, xMSR_IE;
   reg 		   rMSR_BE, xMSR_BE;
   reg 		   ref_rMSR_BIP, xMSR_BIP;
   wire 	   fSKIP = rBRA & !rDLY;
   reg [31:0] 	   rOPA, rOPB;
   always @(rDWBDI or rMXSRC or rPC or rREGA or ref_rRESULT)
     case (rMXSRC)
       2'o0: rOPA <= rREGA;
       2'o1: rOPA <= ref_rRESULT;
       2'o2: rOPA <= rDWBDI;
       2'o3: rOPA <= {rPC, 2'o0};       
     endcase 
   always @(rDWBDI or rMXTGT or rREGB or ref_rRESULT or rSIMM)
     case (rMXTGT)
       2'o0: rOPB <= rREGB;
       2'o1: rOPB <= ref_rRESULT;
       2'o2: rOPB <= rDWBDI;
       2'o3: rOPB <= rSIMM;       
     endcase 
   reg 		    rRES_ADDC;
   reg [31:0] 	    rRES_ADD;
   wire [31:0] 		wADD;
   wire 		wADC;
   wire 		fCCC = !rOPC[5] & rOPC[1]; 
   wire 		fSUB = !rOPC[5] & rOPC[0]; 
   wire 		fCMP = !rOPC[3] & rIMM[1]; 
   wire 		wCMP = (fCMP) ? !wADC : wADD[31]; 
   wire [31:0] 		wOPA = (fSUB) ? ~rOPA : rOPA;
   wire 		wOPC = (fCCC) ? rMSR_C : fSUB;
   assign 		{wADC, wADD} = (rOPB + wOPA) + wOPC; 
   always @(wADC or wADD or wCMP) begin
      {rRES_ADDC, rRES_ADD} <= #1 {wADC, wCMP, wADD[30:0]}; 
   end
   reg [31:0] 	    rRES_LOG;
   always @(rOPA or rOPB or rOPC)
     case (rOPC[1:0])
       2'o0: rRES_LOG <= #1 rOPA | rOPB;
       2'o1: rRES_LOG <= #1 rOPA & rOPB;
       2'o2: rRES_LOG <= #1 rOPA ^ rOPB;
       2'o3: rRES_LOG <= #1 rOPA & ~rOPB;       
     endcase 
   reg [31:0] 	    rRES_SFT;
   reg 		    rRES_SFTC;
   always @(rIMM or rMSR_C or rOPA)
     case (rIMM[6:5])
       2'o0: {rRES_SFT, rRES_SFTC} <= #1 {rOPA[31],rOPA[31:0]};
       2'o1: {rRES_SFT, rRES_SFTC} <= #1 {rMSR_C,rOPA[31:0]};
       2'o2: {rRES_SFT, rRES_SFTC} <= #1 {1'b0,rOPA[31:0]};
       2'o3: {rRES_SFT, rRES_SFTC} <= #1 (rIMM[0]) ? { {(16){rOPA[15]}}, rOPA[15:0], rMSR_C} :
				      { {(24){rOPA[7]}}, rOPA[7:0], rMSR_C};
     endcase 
   wire [31:0] 	    wMSR = {rMSR_C, 3'o0, 
			    20'h0ED32, 
			    4'h0, ref_rMSR_BIP, rMSR_C, ref_rMSR_IE, rMSR_BE};      
   wire 	    fMFSR = (rOPC == 6'o45) & !rIMM[14] & rIMM[0];
   wire 	    fMFPC = (rOPC == 6'o45) & !rIMM[14] & !rIMM[0];
   reg [31:0] 	    rRES_MOV;
   always @(fMFPC or fMFSR or rOPA or rOPB or rPC or rRA
	    or wMSR)
     rRES_MOV <= (fMFSR) ? wMSR :
		 (fMFPC) ? rPC :
		 (rRA[3]) ? rOPB : 
		 rOPA;   
   reg [31:0] 	    rRES_MUL, rRES_MUL0, xRES_MUL;
   always @(rOPA or rOPB) begin
      xRES_MUL <= (rOPA * rOPB);
   end
   always @(posedge gclk)
     if (grst) begin
	rRES_MUL <= 32'h0;
     end else if (rSTALL) begin
	rRES_MUL <= #1 xRES_MUL;	
     end
   reg [31:0] 	 rRES_BSF;
   reg [31:0] 	 xBSRL, xBSRA, xBSLL;
   always @(rOPA or rOPB)
     xBSLL <= rOPA << rOPB[4:0];
   always @(rOPA or rOPB)
     xBSRL <= rOPA >> rOPB[4:0];
   always @(rOPA or rOPB)
     case (rOPB[4:0])
       5'd00: xBSRA <= rOPA;
       5'd01: xBSRA <= {{(1){rOPA[31]}}, rOPA[31:1]};
       5'd02: xBSRA <= {{(2){rOPA[31]}}, rOPA[31:2]};
       5'd03: xBSRA <= {{(3){rOPA[31]}}, rOPA[31:3]};
       5'd04: xBSRA <= {{(4){rOPA[31]}}, rOPA[31:4]};
       5'd05: xBSRA <= {{(5){rOPA[31]}}, rOPA[31:5]};
       5'd06: xBSRA <= {{(6){rOPA[31]}}, rOPA[31:6]};
       5'd07: xBSRA <= {{(7){rOPA[31]}}, rOPA[31:7]};
       5'd08: xBSRA <= {{(8){rOPA[31]}}, rOPA[31:8]};
       5'd09: xBSRA <= {{(9){rOPA[31]}}, rOPA[31:9]};
       5'd10: xBSRA <= {{(10){rOPA[31]}}, rOPA[31:10]};
       5'd11: xBSRA <= {{(11){rOPA[31]}}, rOPA[31:11]};
       5'd12: xBSRA <= {{(12){rOPA[31]}}, rOPA[31:12]};
       5'd13: xBSRA <= {{(13){rOPA[31]}}, rOPA[31:13]};
       5'd14: xBSRA <= {{(14){rOPA[31]}}, rOPA[31:14]};
       5'd15: xBSRA <= {{(15){rOPA[31]}}, rOPA[31:15]};
       5'd16: xBSRA <= {{(16){rOPA[31]}}, rOPA[31:16]};
       5'd17: xBSRA <= {{(17){rOPA[31]}}, rOPA[31:17]};
       5'd18: xBSRA <= {{(18){rOPA[31]}}, rOPA[31:18]};
       5'd19: xBSRA <= {{(19){rOPA[31]}}, rOPA[31:19]};
       5'd20: xBSRA <= {{(20){rOPA[31]}}, rOPA[31:20]};
       5'd21: xBSRA <= {{(21){rOPA[31]}}, rOPA[31:21]};
       5'd22: xBSRA <= {{(22){rOPA[31]}}, rOPA[31:22]};
       5'd23: xBSRA <= {{(23){rOPA[31]}}, rOPA[31:23]};
       5'd24: xBSRA <= {{(24){rOPA[31]}}, rOPA[31:24]};
       5'd25: xBSRA <= {{(25){rOPA[31]}}, rOPA[31:25]};
       5'd26: xBSRA <= {{(26){rOPA[31]}}, rOPA[31:26]};
       5'd27: xBSRA <= {{(27){rOPA[31]}}, rOPA[31:27]};
       5'd28: xBSRA <= {{(28){rOPA[31]}}, rOPA[31:28]};
       5'd29: xBSRA <= {{(29){rOPA[31]}}, rOPA[31:29]};
       5'd30: xBSRA <= {{(30){rOPA[31]}}, rOPA[31:30]};
       5'd31: xBSRA <= {{(31){rOPA[31]}}, rOPA[31]};
     endcase 
   reg [31:0] 	 rBSRL, rBSRA, rBSLL;
   always @(posedge gclk)
     if (grst) begin
	rBSLL <= 32'h0;
	rBSRA <= 32'h0;
	rBSRL <= 32'h0;
     end else if (rSTALL) begin
	rBSRL <= #1 xBSRL;
	rBSRA <= #1 xBSRA;
	rBSLL <= #1 xBSLL;	
     end
   always @(rALT or rBSLL or rBSRA or rBSRL)
     case (rALT[10:9])
       2'd0: rRES_BSF <= rBSRL;
       2'd1: rRES_BSF <= rBSRA;       
       2'd2: rRES_BSF <= rBSLL;
       default: rRES_BSF <= 32'hX;       
     endcase 
   wire 	   fMTS = (rOPC == 6'o45) & rIMM[14] & !fSKIP;
   wire 	   fADDC = ({rOPC[5:4], rOPC[2]} == 3'o0);
   always @(fADDC or fMTS or fSKIP or rMSR_C or rMXALU
	    or rOPA or rRES_ADDC or rRES_SFTC)
     if (fSKIP) begin
	xMSR_C <= rMSR_C;
     end else
       case (rMXALU)
	 3'o0: xMSR_C <= (fADDC) ? rRES_ADDC : rMSR_C;	 
	 3'o1: xMSR_C <= rMSR_C; 
	 3'o2: xMSR_C <= rRES_SFTC; 
	 3'o3: xMSR_C <= (fMTS) ? rOPA[2] : rMSR_C;
	 3'o4: xMSR_C <= rMSR_C;	 
	 3'o5: xMSR_C <= rMSR_C;	 
	 default: xMSR_C <= 1'hX;       
       endcase 
   wire 	    fRTID = (rOPC == 6'o55) & rRD[0] & !fSKIP;   
   wire 	    fRTBD = (rOPC == 6'o55) & rRD[1] & !fSKIP;
   wire 	    fBRK = ((rOPC == 6'o56) | (rOPC == 6'o66)) & (rRA == 5'hC);
   wire 	    fINT = ((rOPC == 6'o56) | (rOPC == 6'o66)) & (rRA == 5'hE);
   always @(fINT or fMTS or fRTID or ref_rMSR_IE or rOPA)
     xMSR_IE <= (fINT) ? 1'b0 :
		(fRTID) ? 1'b1 : 
		(fMTS) ? rOPA[1] :
		ref_rMSR_IE;      
   always @(fBRK or fMTS or fRTBD or ref_rMSR_BIP or rOPA)
     xMSR_BIP <= (fBRK) ? 1'b1 :
		 (fRTBD) ? 1'b0 : 
		 (fMTS) ? rOPA[3] :
		 ref_rMSR_BIP;      
   always @(fMTS or rMSR_BE or rOPA)
     xMSR_BE <= (fMTS) ? rOPA[0] : rMSR_BE;      
   reg [31:0] 	   ref_rRESULT, xRESULT;
   always @(fSKIP or rMXALU or rRES_ADD or rRES_BSF
	    or rRES_LOG or rRES_MOV or rRES_MUL or rRES_SFT)
     if (fSKIP) 
       xRESULT <= 32'h0;
     else
       case (rMXALU)
	 3'o0: xRESULT <= rRES_ADD;
	 3'o1: xRESULT <= rRES_LOG;
	 3'o2: xRESULT <= rRES_SFT;
	 3'o3: xRESULT <= rRES_MOV;
	 3'o4: xRESULT <= (MUL) ? rRES_MUL : 32'hX;	 
	 3'o5: xRESULT <= (BSF) ? rRES_BSF : 32'hX;	 
	 default: xRESULT <= 32'hX;       
       endcase 
   reg [3:0] 	    ref_rDWBSEL, xDWBSEL;
   assign 	    ref_dwb_adr_o = ref_rRESULT[DW-1:2];
   assign 	    ref_dwb_sel_o = ref_rDWBSEL;
   always @(rOPC or wADD)
     case (rOPC[1:0])
       2'o0: case (wADD[1:0]) 
	       2'o0: xDWBSEL <= 4'h8;	       
	       2'o1: xDWBSEL <= 4'h4;	       
	       2'o2: xDWBSEL <= 4'h2;	       
	       2'o3: xDWBSEL <= 4'h1;	       
	     endcase 
       2'o1: xDWBSEL <= (wADD[1]) ? 4'h3 : 4'hC; 
       2'o2: xDWBSEL <= 4'hF; 
       2'o3: xDWBSEL <= 4'h0; 
     endcase 
   reg [14:2] 	    rFSLADR, xFSLADR;   
   assign 	    {ref_fsl_adr_o, ref_fsl_tag_o} = rFSLADR[8:2];
   always @(rALT or rRB) begin
      xFSLADR <= {rALT, rRB[3:2]};      
   end
   always @(posedge gclk)
     if (grst) begin
	ref_rDWBSEL <= 4'h0;
	rFSLADR <= 13'h0;
	rMSR_BE <= 1'h0;
	ref_rMSR_BIP <= 1'h0;
	rMSR_C <= 1'h0;
	ref_rMSR_IE <= 1'h0;
	ref_rRESULT <= 32'h0;
     end else if (gena) begin 
	ref_rRESULT <= #1 xRESULT;
	ref_rDWBSEL <= #1 xDWBSEL;
	rMSR_C <= #1 xMSR_C;
	ref_rMSR_IE <= #1 xMSR_IE;	
	rMSR_BE <= #1 xMSR_BE;	
	ref_rMSR_BIP <= #1 xMSR_BIP;
	rFSLADR <= #1 xFSLADR;
     end
endmodule




module tb;

    // Parameters
    parameter DW = 32;

    // Inputs
    reg [31:0] rREGA, rREGB, rSIMM, rDWBDI;
    reg [1:0] rMXSRC, rMXTGT;
    reg [4:0] rRA, rRB, rRD;
    reg [2:0] rMXALU;
    reg rBRA, rDLY, rSTALL, gclk, grst, gena;
    reg [10:0] rALT;
    reg [15:0] rIMM;
    reg [5:0] rOPC;

    // Outputs
    wire [DW-1:2] ref_dwb_adr_o;
    wire [3:0] ref_dwb_sel_o;
    wire [31:0] ref_rRESULT;
    wire ref_rMSR_IE, ref_rMSR_BIP;

    // Outputs
    wire [DW-1:2] dwb_adr_o;
    wire [3:0] dwb_sel_o;
    wire [31:0] rRESULT;
    wire rMSR_IE, rMSR_BIP;

	wire match;
 	integer total_tests = 0;
	integer failed_tests = 0;

 assign match = (ref_dwb_adr_o === dwb_adr_o) &&  (ref_dwb_sel_o === dwb_sel_o) && (ref_rRESULT === rRESULT) && (ref_rMSR_IE === rMSR_IE) && (ref_rMSR_BIP === rMSR_BIP); 

    // Instantiate the aeMB_xecu module
    ref_aeMB_xecu rf (
        .ref_dwb_adr_o(ref_dwb_adr_o),
        .ref_dwb_sel_o(ref_dwb_sel_o),
        .ref_rRESULT(ref_rRESULT),
        .ref_rMSR_IE(ref_rMSR_IE),
        .ref_rMSR_BIP(ref_rMSR_BIP),
        .rREGA(rREGA),
        .rREGB(rREGB),
        .rMXSRC(rMXSRC),
        .rMXTGT(rMXTGT),
        .rRA(rRA),
        .rRB(rRB),
        .rMXALU(rMXALU),
        .rBRA(rBRA),
        .rDLY(rDLY),
        .rALT(rALT),
        .rSTALL(rSTALL),
        .rSIMM(rSIMM),
        .rIMM(rIMM),
        .rOPC(rOPC),
        .rRD(rRD),
        .rDWBDI(rDWBDI),
        .gclk(gclk),
        .grst(grst),
        .gena(gena)
    );

    // Instantiate the aeMB_xecu module
    aeMB_xecu uut (
        .dwb_adr_o(dwb_adr_o),
        .dwb_sel_o(dwb_sel_o),
        .rRESULT(rRESULT),
        .rMSR_IE(rMSR_IE),
        .rMSR_BIP(rMSR_BIP),
        .rREGA(rREGA),
        .rREGB(rREGB),
        .rMXSRC(rMXSRC),
        .rMXTGT(rMXTGT),
        .rRA(rRA),
        .rRB(rRB),
        .rMXALU(rMXALU),
        .rBRA(rBRA),
        .rDLY(rDLY),
        .rALT(rALT),
        .rSTALL(rSTALL),
        .rSIMM(rSIMM),
        .rIMM(rIMM),
        .rOPC(rOPC),
        .rRD(rRD),
        .rDWBDI(rDWBDI),
        .gclk(gclk),
        .grst(grst),
        .gena(gena)
    );

    // Clock generation
    initial begin
        gclk = 0;
        forever #5 gclk = ~gclk; // 100 MHz clock
    end

    // Test Procedure
    initial begin
        // Initialize inputs
        grst = 1;
        gena = 0;
        rREGA = 0;
        rREGB = 0;
        rMXSRC = 0;
        rMXTGT = 0;
        rRA = 0;
        rRB = 0;
        rMXALU = 0;
        rBRA = 0;
        rDLY = 0;
        rSTALL = 0;
        rSIMM = 0;
        rIMM = 0;
        rOPC = 0;
        rRD = 0;
        rDWBDI = 0;
        rALT = 0;

        // Release reset
        #10 grst = 0;

        // Test Case 1: Simple Addition
        rREGA = 32'h0000000A; // 10
        rREGB = 32'h00000005; // 5
        rMXSRC = 2'b00; // Select rREGA
        rMXTGT = 2'b00; // Select rREGB
        rMXALU = 3'b000; // Add operation
        rOPC = 6'b000000; // ALU operation
        gena = 1;
	compare();
        #10;
        if (rRESULT == 32'h0000000F) begin
            $display("Test Case 1 Passed: Addition Result = %h", rRESULT);
        end else begin
            $display("Test Case 1 Failed: Result = %h", rRESULT);
        end

   repeat (96) begin
      @(posedge gclk);
	rREGA = $random;
	rREGB = $random;
	rSIMM = $random;
	rDWBDI = $random;
	rMXSRC = $random;
	rMXTGT = $random;
	rRA = $random;
	rRB = $random;
	rRD = $random;
	rMXALU = $random;
	rBRA = $random;
	rDLY = $random;
	rSTALL = $random;
	grst = $random;
	gena = $random;
	rALT = $random;
	rIMM = $random;
	rOPC = $random;
     
      compare();
    end
        // Additional test cases can be added similarly...
	$display("All tests passed: design passed");
        $display("\033[1;34mTotal testcases: %d, Failed testcases: %d\033[0m", total_tests, failed_tests);
        // Finish simulation

    if (failed_tests==0) begin
            $display("=====================Your Design Passed======================");
    end
        #100;
        $finish;
    end

task compare;
    begin
        total_tests = total_tests + 1;
        if (match) begin                               //condition to check DUT outputs and calculated //outputs from task are equabegin								
			//$display("\033[1;32mtestcase is passed!!!\033[0m");
			//$display("time = %0t,dwb_adr_o=%h,dwb_sel_o=%h,rRESULT=%h,rMSR_IE=%h,rMSR_BIP=%h\n",$time,dwb_adr_o,dwb_sel_o,rRESULT,rMSR_IE, rMSR_BIP);
			//$display("testcase is passed!!!");
		end

		else begin
			//$display("\033[1;31mtestcase is failed!!!\033[0m");
			//$display("time = %0t,dwb_adr_o=%h,dwb_sel_o=%h,rRESULT=%h,rMSR_IE=%h,rMSR_BIP=%h\n",$time,dwb_adr_o,dwb_sel_o,rRESULT,rMSR_IE, rMSR_BIP);
            failed_tests = failed_tests + 1; 
		end
    end
endtask


    initial begin
        $dumpfile("sim.fsdb");
        $dumpvars(0);
    end

endmodule
